library verilog;
use verilog.vl_types.all;
entity adder_4bit_vlg_vec_tst is
end adder_4bit_vlg_vec_tst;
